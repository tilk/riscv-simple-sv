`ifndef RV_CONFIG
`define RV_CONFIG

import "DPI-C" function string text_mem_file ();
import "DPI-C" function string data_mem_file ();

`endif
